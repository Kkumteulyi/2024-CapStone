module lidar(


	);


/*
UART interface
start cmd : cmd[5] = {0x55, 0xAA, 0x81, 0x00, 0xFA}


*/





